-----------------------------------------------------------------------------------------------------------
-- Floating Point Unit IEEE 754 ( 32 bits support )
-----------------------------------------------------------------------------------------------------------
-- MUX
-- DESCRIPTION : Standard mux
-----------------------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

-----------------------------------------------------------------------------------------------------------

-----------------------------------------------------------------------------------------------------------
-- ENTITY DECLARATION
-----------------------------------------------------------------------------------------------------------

ENTITY MUX IS

    PORT(

        A   :  IN STD_LOGIC; -- INPUT 1
        B   :  IN STD_LOGIC; -- INPUT 2
        Sel :  IN STD_LOGIC; -- SELECTOR
        Z   : OUT STD_LOGIC  -- OUTPUT
    );

END ENTITY;

-----------------------------------------------------------------------------------------------------------

-----------------------------------------------------------------------------------------------------------
-- ARCHITECTURE
-----------------------------------------------------------------------------------------------------------

ARCHITECTURE arch OF MUX IS 


    BEGIN

        Z <= A WHEN Sel = '1' ELSE 
             B;

END ARCHITECTURE;

-----------------------------------------------------------------------------------------------------------