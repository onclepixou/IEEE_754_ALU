-----------------------------------------------------------------------------------------------------------
-- Floating Point Unit IEEE 754 ( 32 bits support )
-----------------------------------------------------------------------------------------------------------
-- Carry look ahead (CLA)
-- DESCRIPTION : sum on 1 bit + carryout
-----------------------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

-----------------------------------------------------------------------------------------------------------

-----------------------------------------------------------------------------------------------------------
-- ENTITY DECLARATION
-----------------------------------------------------------------------------------------------------------

ENTITY CLA IS

    PORT(

        A     :  IN STD_LOGIC; -- Operand 1
        B     :  IN STD_LOGIC; -- Operand 2
        C_IN  :  IN STD_LOGIC; -- IN carry
        C_OUT : OUT STD_LOGIC; -- OUT carry                     
        S     : OUT STD_LOGIC  -- Sum
    );

END ENTITY;

-----------------------------------------------------------------------------------------------------------

-----------------------------------------------------------------------------------------------------------
-- ARCHITECTURE
-----------------------------------------------------------------------------------------------------------

ARCHITECTURE ARCH OF CLA IS 

    SIGNAL c_gen : STD_LOGIC;
    SIGNAL c_pro : STD_LOGIC;
 
    BEGIN

        c_gen <= A AND B;
        c_pro <= A XOR B;

        C_OUT <= c_gen OR ( c_pro AND C_IN );
        S <= c_pro XOR C_IN;

END ARCHITECTURE;

-----------------------------------------------------------------------------------------------------------