-----------------------------------------------------------------------------------------------------------
-- Floating Point Unit IEEE 754 ( 32 bits support )
-----------------------------------------------------------------------------------------------------------
-- COMPUTE BLOCK --> ALU --> ADD_SUB --> ADD_SUB_SIGN_OUT
-- DESCRIPTION : Performs + operation
-----------------------------------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

-----------------------------------------------------------------------------------------------------------

-----------------------------------------------------------------------------------------------------------
-- ENTITY DECLARATION
-----------------------------------------------------------------------------------------------------------

ENTITY ADD_SUB_SIGN_OUT IS

    PORT(

        SA       :  IN STD_LOGIC; -- Augmented operand 1
        SB       :  IN STD_LOGIC; -- Augmented operand 2
        A_BIGGER :  IN STD_LOGIC; -- 1 when A is bigger
        OP_IN    :  IN STD_LOGIC; -- 0 for add, 1 for sub
        OP_OUT   : OUT STD_LOGIC; -- 0 for add, 1 for sub
        SO       : OUT STD_LOGIC  -- Sign out
    );

END ENTITY;

-----------------------------------------------------------------------------------------------------------

-----------------------------------------------------------------------------------------------------------
-- ARCHITECTURE
-----------------------------------------------------------------------------------------------------------

ARCHITECTURE ARCH OF ADD_SUB_SIGN_OUT IS 

    SIGNAL S_AUX : STD_LOGIC;
 
    BEGIN

        S_AUX <= SB XOR OP_IN;

        SO <= SA    WHEN ( A_BIGGER = '1' ) ELSE
              S_AUX WHEN ( A_BIGGER = '0' ) ELSE
              '-';

        OP_OUT <= '1' WHEN SA /= S_AUX else
                  '0';


END ARCHITECTURE;

-----------------------------------------------------------------------------------------------------------